*----------------------------
* NON-INVERTING AMPLIFIER   -
*                           -
* Author: Meel J.           -
* Date: 5 may 2010          -
*----------------------------
*
*--------- NETLISTS ------------------------------*
*
*-- opamp TL084 ----------------------------------*
.inc TL084.cir
Vcc 10 0  DC  15V
Vee 20 0  DC -15V
*       i+ i- V+ V-  O
XTL084   1  0 10 20  21 TL084
*-- amplifier build with TL084 -------------------*
*       i+ i- V+ V-  O
XATL084  1 32 10 20 22 TL084
RF2 22 32 90KOHM
R12 32  0 1KOHM 
*-------------------------------------------------*
*-- opamp TL084 VCVS------------------------------*
.inc opamp84.cir
*       i+ i-  O
Xoa84   1  0  23 opamp84
Rload   23 0  1MEGOhm
*-- amplifier build with TL084 VCVS---------------*
*       i+ i- V+ V-  O
XAoa84  1 34 24 opamp84
RF4 24 34 90KOHM
R14 34  0 1KOHM 
*-------------------------------------------------*
*
*--------- INPUT SOURCE --------------------------*
*
Vin    1 0 AC 1V
*
*--------- ANALYSIS ------------------------------*
*
.AC DEC 100 1HZ 1GHZ
*
*--------- RESULTS -------------------------------*
*
.PROBE
.END