* Z:\home\dries\Projects\SignaalVerwerking\ideaal.ascz
R3 N006 vin 19894
R1 N002 N005 19894
R2 N004 N003 19894
C2 Vout N004 1n
C1 N003 N002 21.33n
R6 N005 N001 19894
R4 N003 N006 19894
R5 Vout N001 59683
V1 vin 0 AC 1
XU4 N001 N006 N005 opampIdeal
XU5 N002 0 N003 opampIdeal
XU6 N004 0 Vout opampIdeal
.ac dec 100 100 1MEG
.lib Z:\home\dries\Projects\SignaalVerwerking\docs\OpampModel\OPAMP_PSPICE\opampIdeal.cir
.backanno
.end
