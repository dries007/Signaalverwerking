* Bode (LTSpice export)
.inc opampIdeaal.cir

.model r res(r = 1 DEV 1%)
.model c cap(c = 1 DEV 1%)

R1 N001 vin r 6.1426K
V1 vin 0 AC 1
XU1 N001 0 N002 opampIdeal
C1 N002 N001 c 1e-8
R2 N002 N001 r 26.648K
R3 vout N001 r 8.6869K
XU2 N003 0 N004 opampIdeal
XU3 N005 0 vout opampIdeal
R4 N003 N002 r 8.6869K
R5 N005 N004 r 8.6869K
R6 vout N005 r 8.6869K
C2 N004 N003 c 1e-8

.ac dec 100 100 1MEG
.mc 10 AC V(R6) YMAX LIST OUTPUT ALL
.probe
.end
