* Z:\home\dries\Projects\SignaalVerwerking\vcvs.asc
R3 N006 vin 19894
R1 N002 N005 19894
R2 N004 N003 19894
C2 Vout N004 1n
C1 N003 N002 21.33n
R6 N005 N001 19894
R4 N003 N006 19894
R5 Vout N001 59683
V1 vin 0 AC 1
XU1 N001 N006 N005 opamp84
XU2 N002 0 N003 opamp84
XU3 N004 0 Vout opamp84
.ac dec 100 100 1MEG
.lib Z:\home\dries\Projects\SignaalVerwerking\docs\OpampModel\OPAMP_PSPICE\opamp84.cir
.backanno
.end
