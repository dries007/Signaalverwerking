* H ideaal
.inc tl084.cir
.model rmod res(r = 1 DEV/GAUSS 1%)
.model cmod cap(c = 1 DEV/GAUSS 1%)
R3 6 vin rmod 19894
R1 2 5 rmod 19894
R2 4 3 rmod 19894
C2 Vout 4 cmod 1n
C1 3 2 cmod 21.33n
R6 5 1 rmod 19894
R4 3 6 rmod 19894
R5 Vout 1 rmod 59683
V1 vin 0 AC 1
V2 vp 0 15
V3 0 vn 15
XU4 1 6 vp vn 5 tl084
XU5 2 0 vp vn 3 tl084
XU6 4 0 vp vn Vout tl084
.ac dec 100 100 1MEG
.mc 10 ac V(V1) ymax list output all
.probe					  
.end
